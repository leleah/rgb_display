module main(
input Clock,
output reg [4:0] Red,
output reg  [5:0] Green,
output reg  [4:0] Blue,
output reg  Vsync,
output reg  Hsync,
output reg  Pixel_Clock,
output reg  DEN
);

always @(posedge Clock) begin


end

endmodule
